/*  written by      :   Mohamed S. Helal
    date created   	:   Mar, 9th, 2025
    description     :   FFT input ROM, reads a file "testvecROM.txt"
                        containing 64 decimal numbers.
	>>important		:	it reads reverse bit order for the first 3 bits
    version         :   0.0
*/

module FFT_xn_ROM (
    input   wire        clk,
    input   wire [5:0]  addr,   // 6-bit address (since 2^6 = 64)
    output  reg  [15:0] dout    // 16-bit output
);

// Internal memory array to store 64 values
reg [15:0] rom [0:63];

// File read operation
initial begin
    $readmemh("testvecROM.txt", rom);  // Read signed hex numbers (generated by Octave)
end

// Read operation
always @(*) begin
    dout = rom[{addr[5:3],addr[0],addr[1],addr[2]}];	// read 0>4>2>6>1>5>3>7>8>12...etc
end

endmodule
